AND gates

.include  ..\gpdk90nm\gpdk90nm_tt.cir

.subckt 2inAND in1 in2 out1 Vdd Vss Len Ratio

.end

.subckt 3inAND in1 in2 in3 out1 Vdd Vss Len Ratio

.end
