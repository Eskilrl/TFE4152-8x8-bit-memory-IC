*Bitcell

.include logic_gates_library.cir

*Parameters

.param Vdd=0.3V

.param L1=1u
.param W1=10u

.subckt SRlatch inp outp Vdd Vss
xNAND1 inp !Q Q Vdd Vss 2inNAND
xNOT1 inp !inp Vdd Vss 1inNOT
xNAND2 Q !inp !Q Vdd Vss 2inNAND
.ends

*Test

V1 1 0 dc Vdd
Vin in 0 dc 0 

xAND1 in 1 Y 1 0 2inAND

.dc Vin 0 Vdd 0.01
.plot v(Y)
