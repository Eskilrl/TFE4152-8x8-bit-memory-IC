module FlipFlop (

//Inputs

input i_sel,
input i_inp,
input i_wr,

//OUPUTS

ouptut o_outp
);







endmodule
