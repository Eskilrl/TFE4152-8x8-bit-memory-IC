*Bitcell

.include logic_gates_library.cir

*Parameters

.param Vdd=1

.param L1=1u
.param W1=10u

.subckt SRlatch inp notoutp Vdd Vss
xNOR1 inp notoutp outp Vdd Vss 2inNOR
xNOT1 inp notinp Vdd Vss 1inNOT
xNOR2 outp notinp notoutp Vdd Vss 2inNOR
.ends

.subckt SRbitcell inp sel rw outp Vdd Vss
xAND1 inp sel rw tempinp Vdd Vss 3inAND
xNOT1 rw notrw Vdd Vss 1inNOT
xSR1 tempinp tempoutp Vdd Vss SRlatch
xAND2 tempoutp notrw sel outp Vdd Vss 3inAND
.ends

*Test

V1 1 0 dc Vdd
Vinp inp 0 PULSE(0 Vdd 15ns 0.1ns 0.1ns 10ns 30ns)
*Vsel sel 0 PULSE(0 Vdd 9ns 0.1ns 0.1ns 2ns 15ns)
*Vrw rw 0 PULSE(0 Vdd 10ns 0.1ns 0.1ns 10ns 20ns)

xSR1 inp Y 1 0 SRlatch
*xBitcell inp sel rw Y 1 0 SRbitcell

.tran 5n 40n
.plot v(inp) v(Y)



